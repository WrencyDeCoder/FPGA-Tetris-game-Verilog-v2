module score_digit_rom (
    input  wire [3:0]  number,     // 0–9
    output wire [79:0] data        // 10  * 8 
);

    // 10 digit * 80 bit/digit = 800 bit
    localparam [800-1:0] ROM = {
        //======================
        // 9
        //======================
            8'b01111100, 8'b11000110, 8'b11000110, 8'b11000110,
            8'b01111110, 8'b00000110, 8'b00000110, 8'b00001100,
            8'b00011000, 8'b01110000,
				
        //======================
        // 8
        //======================
            8'b01111100, 8'b11000110, 8'b11000110, 8'b01111100,
            8'b11000110, 8'b11000110, 8'b11000110, 8'b11000110,
            8'b11000110, 8'b01111100,
       
        //======================
        // 7
        //======================
            8'b11111110, 8'b11000110, 8'b00000110, 8'b00001100,
            8'b00011000, 8'b00110000, 8'b01100000, 8'b01100000,
            8'b01100000, 8'b01100000,

        //======================
        // 6
        //======================
            8'b00111000, 8'b01100000, 8'b11000000, 8'b11111100,
            8'b11000110, 8'b11000110, 8'b11000110, 8'b11000110,
            8'b11000110, 8'b01111100,
       
        //======================
        // 5
        //======================
            8'b11111110, 8'b11000000, 8'b11000000, 8'b11111100,
            8'b00000110, 8'b00000110, 8'b00000110, 8'b11000110,
            8'b11000110, 8'b01111100,

        //======================
        // 4
        //======================
            8'b00001100, 8'b00011100, 8'b00111100, 8'b01101100,
            8'b11001100, 8'b11111110, 8'b00001100, 8'b00001100,
            8'b00001100, 8'b00001100,
       
        //======================
        // 3
        //======================
            8'b01111100, 8'b11000110, 8'b00000110, 8'b00001100,
            8'b00111100, 8'b00001100, 8'b00000110, 8'b00000110,
            8'b11000110, 8'b01111100,
    
        //======================
        // 2
        //======================
            8'b01111100, 8'b11000110, 8'b00000110, 8'b00001100,
            8'b00011000, 8'b00110000, 8'b01100000, 8'b11000000,
            8'b11000110, 8'b11111110,
  
        //======================
        // 1
        //======================
            8'b00011000, 8'b00111000, 8'b01111000, 8'b00011000,
            8'b00011000, 8'b00011000, 8'b00011000, 8'b00011000,
            8'b00011000, 8'b01111110,
      
        //======================
        // 0
        //======================
            8'b01111100, 8'b11000110, 8'b11001110, 8'b11011110,
            8'b11110110, 8'b11100110, 8'b11000110, 8'b11000110,
            8'b11000110, 8'b01111100
    };

    // access digit
    assign data = ROM[number*80 +: 80];

endmodule
