//======================================================
// game_over_text_rom.v
//======================================================
module game_over_text_rom (
    input  wire [9:0] X,
    input  wire [9:0] Y,

    output wire inside_area,
    output reg  is_pixel
);

    localparam integer TEXT_W = 166;
    localparam integer TEXT_H = 16;

    localparam integer MSG_X = 30;
    localparam integer MSG_Y = 180;

    // 166-bit per row (6 + 32*5)
    reg [TEXT_W-1:0] text_bitmap [0:TEXT_H-1];

    initial begin

        // ---------------- ROW 0 ----------------
        text_bitmap[0] = {
            6'b001111,
            32'b11111111111111000111111111111110,
            32'b00111111000000001111111000111111,
            32'b11111111100000000000000011111111,
            32'b11111100011111100000111111100011,
            32'b11111111111111011111111111111110
        };

        // ---------------- ROW 1 ----------------
        text_bitmap[1] = {
            6'b011111,
            32'b11111111110011111111111111100011,
            32'b11111000000000111111100111111111,
            32'b11111111000000000000000111111111,
            32'b11111100011111100000111111100111,
            32'b11111111111111011111111111111110
        };

        // ---------------- ROW 2 ----------------
        text_bitmap[2] = {
            6'b111111,
            32'b11111110111111111111111110000111,
            32'b11111011111111111111111100000000,
            32'b00001111111111111011111110000011,
            32'b11111011111111111111011111111111,
            32'b0111111111111111110
        };

        // ---------------- ROW 3 ----------------
        text_bitmap[3] = {
            6'b111111,
            32'b00000000000111111000001111111011,
            32'b11111111011111111110111111000000,
            32'b00000000000000111111000001111111,
            32'b01111110000011111110111111000000,
            32'b00000001111110000011111110
        };

        // ---------------- ROW 4 ----------------
        text_bitmap[4] = {
            6'b111111,
            32'b00000000000111111000001111111011,
            32'b11111111011111111110111111000000,
            32'b00000000000000111111000001111111,
            32'b01111110000011111110111111000000,
            32'b00000001111110000011111110
        };

        // ---------------- ROW 5 ----------------
        text_bitmap[5] = {
            6'b111111,
            32'b00000000000111111000001111111011,
            32'b11111111111111111110111111000000,
            32'b00000000000000111111000001111111,
            32'b01111110000011111110111111000000,
            32'b00000001111110000011111110
        };

        // ---------------- ROW 6 ----------------
        text_bitmap[6] = {
            6'b111111,
            32'b00000000000111111000001111111011,
            32'b11111111111111111110111111000000,
            32'b00000000000000111111000001111111,
            32'b01111110000011111110111111000000,
            32'b00000001111110000011111110
        };

        // ---------------- ROW 7 ----------------
        text_bitmap[7] = {
            6'b111111,
            32'b00111111100011111111111111101111,
            32'b11111111110111111111110000000000,
            32'b00000000111111000001111111011111,
            32'b10000011111110111111111110000000,
            32'b0111111111111111000
        };

        // ---------------- ROW 8 ----------------
        text_bitmap[8] = {
            6'b111111,
            32'b00111111100011111111111111101111,
            32'b11001111101111111111100000000000,
            32'b00000000111111000001111111011111,
            32'b10000111111110111111111110000000,
            32'b0111111111111111000
        };

        // ---------------- ROW 9 ----------------
        text_bitmap[9] = {
            6'b111111,
            32'b00111111111011111111111111101111,
            32'b11000010001111111111100000000000,
            32'b00000000111111000001111111001111,
            32'b11000011111111001111111111000000,
            32'b0111111111111111000
        };

        // ---------------- ROW 10 ----------------
        text_bitmap[10] = {
            6'b111111,
            32'b00000111111011111100000111111011,
            32'b11110000100011111100000000000000,
            32'b00000000111111000001111111011111,
            32'b10001111111100001111110000000000,
            32'b01111110000011111110
        };

        // ---------------- ROW 11 ----------------
        text_bitmap[11] = {
            6'b111111,
            32'b00000111111011111100000111111011,
            32'b11110000000011111100000000000000,
            32'b00000000111111000001111111111111,
            32'b00001111110000000000111111000000,
            32'b01111110000011111110
        };

        // ---------------- ROW 12 ----------------
        text_bitmap[12] = {
            6'b111111,
            32'b00000111111011111100000111111011,
            32'b11110000000011111100000000000000,
            32'b00000000111111000001111111111110,
            32'b00001111110000000000111111000000,
            32'b01111110000011111110
        };

        // ---------------- ROW 13 ----------------
        text_bitmap[13] = {
            6'b111111,
            32'b11111111011111110000011111101111,
            32'b11000000001111111011111111100000,
            32'b00000000111111111111111011111111,
            32'b10000001111111111111111011111100,
            32'b00001111110000011111110
        };

        // ---------------- ROW 14 ----------------
        text_bitmap[14] = {
            6'b011111,
            32'b11111110001111110000011111101111,
            32'b11000000001111111001111111110000,
            32'b00000000111111111111110001111111,
            32'b10000000011111111111111011111100,
            32'b00001111110000011111110
        };

        // ---------------- ROW 15 ----------------
        text_bitmap[15] = {
            6'b001111,
            32'b11111110001111110000011111101111,
            32'b11000000001111111000111111110000,
            32'b00000000111111111111100001111111,
            32'b10000000001111111111111011111100,
            32'b00001111110000011111110
        };
    end

    // -------------------------------------------
    // Inside display area
    // -------------------------------------------
    assign inside_area =
        (X >= MSG_X) && (X < MSG_X + TEXT_W) &&
        (Y >= MSG_Y) && (Y < MSG_Y + TEXT_H);

    // -------------------------------------------
    // Pixel fetch
    // -------------------------------------------
    always @(*) begin
        if (inside_area)
            is_pixel = text_bitmap[Y - MSG_Y][TEXT_W - 1 - (X - MSG_X)];
        else
            is_pixel = 1'b0;
    end

endmodule
